`ifndef FIFO_IN_SEQUENCER_SV
`define FIFO_IN_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(fifo_in_tx) fifo_in_sequencer_t;


`endif // FIFO_IN_SEQUENCER_SV
