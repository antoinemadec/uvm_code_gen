`ifndef AHB_SEQUENCER_SV
`define AHB_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(ahb_tx) ahb_sequencer_t;


`endif // AHB_SEQUENCER_SV
