`ifndef HANDSHAKE_SEQUENCER_SV
`define HANDSHAKE_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(handshake_tx) handshake_sequencer_t;


`endif // HANDSHAKE_SEQUENCER_SV
