package ahb_pkg;

  `include "uvm_macros.svh"

  import uvm_pkg::*;


  `include "ahb_tx.sv"
  `include "ahb_config.sv"
  `include "ahb_driver.sv"
  `include "ahb_monitor.sv"
  `include "ahb_sequencer.sv"
  `include "ahb_coverage.sv"
  `include "ahb_agent.sv"
  `include "ahb_seq_lib.sv"

endpackage : ahb_pkg
